-- Processador Versao: 04/11/2024

libraRY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cpu is
	port( 
			clk			: in	std_LOGIC;
			reset			: in	std_LOGIC;
			wait2			: in	std_LOGIC;
			entrada     : in  std_logic_vector(7 downto 0);
			saidaREAL   : out std_logic_vector(7 downto 0);
			saidaRR     : out std_logic_vector(7 downto 0);
			saidaA      : out std_logic_vector(7 downto 0);
			zero			: out	std_LOGIC;
			maior			: out	std_LOGIC;
			menor			: out	std_LOGIC;
			LED1			: out	std_LOGIC := '0';
			LED2			: out	std_LOGIC := '0';
			LED3			: out	std_LOGIC := '0';
			LED4			: out	std_LOGIC := '0';
			LED5			: out	std_LOGIC := '0';
			over			: out	std_LOGIC
		);
end cpu;

ARCHITECTURE main of cpu is

	TYPE STATES				is (fetch, fetch2, decode, exec, exec2);						-- Estados da Maquina de Controle do Processador
	
	signal RA : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal RB : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal RR : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal PC : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal IR : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	
	CONSTANT ADD       : STD_LOGIC_VECTOR(3 downto 0) := "0000";
	CONSTANT SUB       : STD_LOGIC_VECTOR(3 downto 0) := "0001";
	CONSTANT AND1      : STD_LOGIC_VECTOR(3 downto 0) := "0010";
	CONSTANT OR1       : STD_LOGIC_VECTOR(3 downto 0) := "0011";
	CONSTANT NOT1      : STD_LOGIC_VECTOR(3 downto 0) := "0100";
	CONSTANT CMP       : STD_LOGIC_VECTOR(3 downto 0) := "0101";
	CONSTANT JMP       : STD_LOGIC_VECTOR(3 downto 0) := "0110";
	CONSTANT JEQ       : STD_LOGIC_VECTOR(3 downto 0) := "0111";
	CONSTANT JGR       : STD_LOGIC_VECTOR(3 downto 0) := "1000";
	CONSTANT LOAD      : STD_LOGIC_VECTOR(3 downto 0) := "1001";
	CONSTANT STORE     : STD_LOGIC_VECTOR(3 downto 0) := "1010";
	CONSTANT MOV       : STD_LOGIC_VECTOR(3 downto 0) := "1011";
	CONSTANT IN1       : STD_LOGIC_VECTOR(3 downto 0) := "1100";
	CONSTANT OUT1      : STD_LOGIC_VECTOR(3 downto 0) := "1101";
	CONSTANT WAIT1     : STD_LOGIC_VECTOR(3 downto 0) := "1110";
	CONSTANT MY        : STD_LOGIC_VECTOR(3 downto 0) := "1111";
	
	signal ESPERA : STD_LOGIC := '0';
	
	signal X : STD_LOGIC_VECTOR (7 downto 0) := (others => '0'); --Operadores da ULA
	signal Y : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal RESULT   : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
	signal INIT_ULA : STD_LOGIC := '0';
	signal FRzero   : STD_LOGIC := '0';
	signal FRmaior  : STD_LOGIC := '0';
	signal FRmenor  : STD_LOGIC := '0';
	signal FRover   : STD_LOGIC := '0';
	                  
	signal data_in    : std_logic_vector(7 downto 0) := (others => '0');
	signal raddress   : std_logic_vector(7 downto 0) := (others => '0');
	signal waddress   : std_logic_vector(7 downto 0) := (others => '0');
	signal write1     : std_logic := '0';                   
	signal data_out   : std_logic_vector(7 downto 0) := (others => '0');
	
	component ram256x8
			port(
				clock		: IN STD_LOGIC  := '1';
				data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
				rdaddress		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
				wraddress		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
				wren		: IN STD_LOGIC  := '0';
				q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
			);
	end component;


begin
	    ram_instance: ram256x8
        port map (
            clock     => (NOT clk),
            data      => data_in,      
            rdaddress => raddress,     
            wraddress => waddress,     
            wren      => write1,     
            q         => data_out
        );

-- Maquina de Controle
process(clk, reset)

	variable state : STATES := fetch;

begin

IF(reset = '1') THEN

	RA <= (others => '0');
	RB <= (others => '0');
	RR <= (others => '0');
	PC <= (others => '0');
	IR <= (others => '0');
	saidaREAL <= (others => '0');

	data_in  <= (others => '0');
	waddress <= (others => '0');
	write1   <= '0';
	state := fetch;
	
	LED1	<= '0';
	LED2	<= '0';
	LED3	<= '0';
	LED4	<= '0';
	LED5	<= '0';

ELSIF(rising_edge(clk)) THEN
		
		IF(INIT_ULA = '1') THEN --Controle das saidas da ULA
			RR <= RESULT;
			INIT_ULA <= '0';
		END IF;	
			
		case state is
		
--************************************************************************
-- FETCH STATE
--************************************************************************		
		
		when fetch =>
		
		LED1	<= '1';
		LED2	<= '0';
		LED3	<= '0';
		LED4	<= '0';
		LED5	<= '0';
		
			-- Inicio das acoes do ciclo de Busca !!       
			raddress <= PC;
			STATE := fetch2;
			
-- XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX

--************************************************************************
-- FETCH2 STATE
--************************************************************************		
		
		when fetch2 =>
		
		LED1	<= '0';
		LED2	<= '1';
		LED3	<= '0';
		LED4	<= '0';
		LED5	<= '0';
		
			-- Inicio das acoes do ciclo de Busca !!       
			IR <= data_out;
			--saidaA <= data_out;
			saidaREAL <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
			PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

			STATE := decode;
			
-- XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX  
        			

--************************************************************************
-- DECODE STATE
--************************************************************************
		when decode =>
		
		LED1	<= '0';
		LED2	<= '0';
		LED3	<= '1';
		LED4	<= '0';
		LED5	<= '0';

--========================================================================
-- ADD ou SUB ou AND ou OR ou CMP
--========================================================================			
			IF(IR(7 DOWNTO 4) = ADD or (IR(7 DOWNTO 4) = "0001") or (IR(7 DOWNTO 4) = "0010")
				 or (IR(7 DOWNTO 4) = "0011") or (IR(7 DOWNTO 4) = "0101")) THEN
				 
				 IF((IR(3 DOWNTO 0) = "0000")) THEN  -- A A
					  X <= RA;
					  Y <= RA;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "0001") THEN  -- A B
					  X <= RA;
					  Y <= RB;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "0011") THEN  -- A i
					  X <= RA;
					  raddress <= PC;
				 ELSIF(IR(3 DOWNTO 0) = "0010") THEN  -- A R
					  X <= RA;
					  Y <= RR;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "0100") THEN  -- B A
					  X <= RB;
					  Y <= RA;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "0101") THEN  -- B B
					  X <= RB;
					  Y <= RB;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "0111") THEN  -- B i
					  X <= RB;
					  raddress <= PC;
				 ELSIF(IR(3 DOWNTO 0) = "0110") THEN  -- B R
					  X <= RB;
					  Y <= RR;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "1100") THEN  -- i A
					  raddress <= PC;
					  Y <= RA;
				 ELSIF(IR(3 DOWNTO 0) = "1101") THEN  -- i B
					  raddress <= PC;
					  Y <= RB;
				 ELSIF(IR(3 DOWNTO 0) = "1110") THEN  -- i R
					  raddress <= PC;
					  Y <= RR;
				 ELSIF(IR(3 DOWNTO 0) = "1000") THEN  -- R A
					  X <= RR;
					  Y <= RA;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "1001") THEN  -- R B
					  X <= RR;
					  Y <= RB;
					  INIT_ULA <= '1';
				 ELSIF(IR(3 DOWNTO 0) = "1011") THEN  -- R i
					  X <= RR;
					  raddress <= PC;
				 ELSIF(IR(3 DOWNTO 0) = "1010") THEN  -- R R
					  X <= RR;
					  Y <= RR;
					  INIT_ULA <= '1';
				 END IF;
				 state := exec;
			END IF;

--========================================================================
-- NOT
--========================================================================			
			IF(IR(7 DOWNTO 4) = NOT1) THEN
				IF(IR(3 DOWNTO 2) = "00") THEN
					X <= RA;
					INIT_ULA <= '1';
				ELSIF(IR(3 DOWNTO 2) = "01") THEN
					X <= RB;
					INIT_ULA <= '1';
				ELSIF(IR(3 DOWNTO 2) = "10") THEN
					X <= RR;
					INIT_ULA <= '1';
				ELSIF(IR(3 DOWNTO 2) = "11") THEN
					raddress <= PC;
				END IF;
				
				state := exec;
			END IF;

--========================================================================
-- JMP
--========================================================================		
			IF(IR(7 DOWNTO 4) = JMP) THEN
				raddress <= PC;
				state := exec;
			END IF;
			
--========================================================================
-- JEQ
--========================================================================			
			IF(IR(7 DOWNTO 4) = JEQ) THEN
				IF(FRzero = '1') THEN
					raddress <= PC;
				END IF;
				state := exec;
			END IF;
			

--========================================================================
-- JGR
--========================================================================			
			IF(IR(7 DOWNTO 4) = JGR) THEN
				IF(FRzero = '0' and FRmaior ='1') THEN
					raddress <= PC;
				END IF;
				state := exec;
			END IF;
			
--========================================================================
-- LOAD
--========================================================================            
			IF (IR(7 DOWNTO 4) = LOAD) THEN

				 IF (IR(3 DOWNTO 0) = "0000") THEN  -- A A: Carrega para o registrador RA o conteúdo do endereço em RA
					  raddress <= RA;

				 ELSIF (IR(3 DOWNTO 0) = "0001") THEN  -- A B: Carrega para o registrador RA o conteúdo do endereço em RB
					  raddress <= RB;

				 ELSIF (IR(3 DOWNTO 0) = "0011") THEN  -- A i: Carrega para o registrador RA o conteúdo do endereço imediato
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "0010") THEN  -- A R: Carrega para o registrador RA o valor do endereço em RR
					  raddress <= RR;

				 ELSIF (IR(3 DOWNTO 0) = "0100") THEN  -- B A: Carrega para o registrador RB o conteúdo do endereço em RA
					  raddress <= RA;

				 ELSIF (IR(3 DOWNTO 0) = "0101") THEN  -- B B: Carrega para o registrador RB o conteúdo do endereço em RB
					  raddress <= RB;

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i: Carrega para o registrador RB o conteúdo do endereço imediato
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "0110") THEN  -- B R: Carrega para o registrador RB o valor do endereço em RR
					  raddress <= RR;

				 ELSIF (IR(3 DOWNTO 0) = "1000") THEN  -- R A: Carrega para o registrador RR o conteúdo do endereço em RA
					  raddress <= RA;

				 ELSIF (IR(3 DOWNTO 0) = "1001") THEN  -- R B: Carrega para o registrador RR o conteúdo do endereço em RB
					  raddress <= RB;

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i: Carrega para o registrador RR o conteúdo do endereço imediato
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "1010") THEN  -- R R: Carrega para o registrador RR o valor do endereço em RR
					  raddress <= RR;

				 END IF;
				 state := exec;
			END IF;

--========================================================================
-- STORE
--========================================================================            
			IF (IR(7 DOWNTO 4) = STORE) THEN

				 IF (IR(3 DOWNTO 0) = "0000") THEN  -- A A: 
					  waddress <= RA;
					  data_in <= RA;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0001") THEN  -- A B: 
					  waddress <= RB;
					  data_in <= RA;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0010") THEN  -- A R:
					  waddress <= RR;
					  data_in <= RA;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0011") THEN  -- A i:
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "0100") THEN  -- B A: 
					  waddress <= RA;
					  data_in <= RB;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0101") THEN  -- B B: 
					  waddress <= RB;
					  data_in <= RB;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0110") THEN  -- B R:
					  waddress <= RR;
					  data_in <= RB;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i:
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "1000") THEN  -- R A:
					  waddress <= RA;
					  data_in <= RR;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "1001") THEN  -- R B:
					  waddress <= RB;
					  data_in <= RR;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "1010") THEN  -- R R:
					  waddress <= RR;
					  data_in <= RR;
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i:
					  raddress <= PC;

				 END IF;

				 state := exec;

			END IF;

			

--========================================================================
-- MOV
--========================================================================         
			IF (IR(7 DOWNTO 4) = MOV) THEN

				 IF (IR(3 DOWNTO 0) = "0001") THEN  -- A B: Move o valor de RB para RA
					  RA <= RB;

				 ELSIF (IR(3 DOWNTO 0) = "0010") THEN  -- A R: Move o valor de RR para RA
					  RA <= RR;

				 ELSIF (IR(3 DOWNTO 0) = "0011") THEN  -- A i: Move o valor imediato para RA
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "0100") THEN  -- B A: Move o valor de RA para RB
					  RB <= RA;

				 ELSIF (IR(3 DOWNTO 0) = "0110") THEN  -- B R: Move o valor de RR para RB
					  RB <= RR;

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i: Move o valor imediato para RB
					  raddress <= PC;

				 ELSIF (IR(3 DOWNTO 0) = "1000") THEN  -- R A: Move o valor de RA para RR
					  RR <= RA;

				 ELSIF (IR(3 DOWNTO 0) = "1001") THEN  -- R B: Move o valor de RB para RR
					  RR <= RB;

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i: Move o valor imediato para RR
					  raddress <= PC;
				 END IF;

				 state := exec;
			END IF;
			
--========================================================================
-- IN
--========================================================================            
			IF (IR(7 DOWNTO 4) = IN1) THEN

				 IF (IR(3 DOWNTO 2) = "00") THEN  -- A
					  RA <= entrada;

				 ELSIF (IR(3 DOWNTO 2) = "01") THEN  -- B
					  RB <= entrada;

				 ELSIF (IR(3 DOWNTO 2) = "10") THEN  -- R
					  RR <= entrada;

				 END IF;
					state := fetch;
			END IF;
			
--========================================================================
-- OUT
--========================================================================            
			IF (IR(7 DOWNTO 4) = OUT1) THEN

				 IF (IR(3 DOWNTO 2) = "00") THEN  -- A
					  saidaREAL <= RA;

				 ELSIF (IR(3 DOWNTO 2) = "01") THEN  -- B
					  saidaREAL <= RB;

				 ELSIF (IR(3 DOWNTO 2) = "10") THEN  -- R
					  saidaREAL <= RR;

				 END IF;
					state := fetch;
			END IF;

--========================================================================
-- WAIT
--========================================================================            
			IF (IR(7 DOWNTO 4) = WAIT1) THEN
				IF(ESPERA = '0') THEN
					ESPERA <= '1';
					state := decode;
				ELSE
					IF(WAIT2 = '1') THEN
						ESPERA <= '0';
						state := fetch;
					END IF;
				END IF;
			END IF;

-- XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX		

					
							
		
								
							
								

--************************************************************************
-- EXECUTE STATE
--************************************************************************								
					
			when exec =>
			
			LED1	<= '0';
			LED2	<= '0';
			LED3	<= '0';
			LED4	<= '1';
			LED5	<= '0';

--========================================================================
-- EXEC ADD ou SUB ou AND ou OR ou CMP
--========================================================================			
			IF (IR(7 DOWNTO 4) = ADD OR (IR(7 DOWNTO 4) = "0001") OR (IR(7 DOWNTO 4) = "0010") OR 
				 (IR(7 DOWNTO 4) = "0011") OR (IR(7 DOWNTO 4) = "0101")) THEN

				 IF (IR(3 DOWNTO 0) = "0011") THEN  -- A i
					  Y <= data_out;
					  --RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  INIT_ULA <= '1';
					  
				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i
					  Y <= data_out;
					  --RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  INIT_ULA <= '1';
					  
				 ELSIF (IR(3 DOWNTO 0) = "1100") THEN  -- i A
					  X <= data_out;
					  --RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  INIT_ULA <= '1';
					  
				 ELSIF (IR(3 DOWNTO 0) = "1101") THEN  -- i B
					  X <= data_out;
					  --RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  INIT_ULA <= '1';
					  
				 ELSIF (IR(3 DOWNTO 0) = "1110") THEN  -- i R
					  Y <= data_out;
					  --RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  INIT_ULA <= '1';
					  
				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i
					  Y <= data_out;
					  --RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  INIT_ULA <= '1';
					  
				 END IF;

				 state := fetch;

			END IF;

--========================================================================
-- NOT
--========================================================================			
			IF(IR(7 DOWNTO 4) = NOT1) THEN
				IF(IR(3 DOWNTO 2) = "11") THEN
					X <= data_out;
					PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					INIT_ULA <= '1';
				END IF;
				
				state := fetch;
			END IF;
			
--========================================================================
-- JMP
--========================================================================		
			IF(IR(7 DOWNTO 4) = JMP) THEN
				PC <= data_out;
				state := fetch;
			END IF;

--========================================================================
-- JEQ
--========================================================================			
			IF(IR(7 DOWNTO 4) = JEQ) THEN
				IF(FRzero = '1') THEN
					PC <= data_out;
				ELSE
					PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
				END IF;
				state := fetch;
			END IF;
			
--========================================================================
-- JGR
--========================================================================			
			IF(IR(7 DOWNTO 4) = JGR) THEN
				IF(FRzero = '0' and FRmaior ='1') THEN
					PC <= data_out;
				ELSE
					PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
				END IF;
				state := fetch;
			END IF;
			
--========================================================================
-- LOAD
--========================================================================            
			IF (IR(7 DOWNTO 4) = LOAD) THEN

				 IF (IR(3 DOWNTO 0) = "0000") THEN  -- A A: Carrega para o registrador RA o conteúdo do endereço em RA
					  RA <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "0001") THEN  -- A B: Carrega para o registrador RA o conteúdo do endereço em RB
					  RA <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "0011") THEN  -- A i: Carrega para o registrador RA o valor imediato
					  raddress <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

				 ELSIF (IR(3 DOWNTO 0) = "0010") THEN  -- A R: Carrega para o registrador RA o conteúdo do endereço em RR
					  RA <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "0100") THEN  -- B A: Carrega para o registrador RB o conteúdo do endereço em RA
					  RB <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "0101") THEN  -- B B: Carrega para o registrador RB o conteúdo do endereço em RB
					  RB <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i: Carrega para o registrador RB o valor imediato
					  raddress <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

				 ELSIF (IR(3 DOWNTO 0) = "0110") THEN  -- B R: Carrega para o registrador RB o conteúdo do endereço em RR
					  RB <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "1000") THEN  -- R A: Carrega para o registrador RR o conteúdo do endereço em RA
					  RR <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "1001") THEN  -- R B: Carrega para o registrador RR o conteúdo do endereço em RB
					  RR <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i: Carrega para o registrador RR o valor imediato
					  raddress <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

				 ELSIF (IR(3 DOWNTO 0) = "1010") THEN  -- R R: Carrega para o registrador RR o conteúdo do endereço em RR
					  RR <= data_out;

				 END IF;
				 state := exec2;
			END IF;
		
--========================================================================
-- STORE
--========================================================================            
			IF (IR(7 DOWNTO 4) = STORE) THEN
				 

				 IF (IR(3 DOWNTO 0) = "0011") THEN  -- A i:
					  waddress <= data_out;
					  data_in <= RA;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i:
					  waddress <= data_out;
					  data_in <= RB;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  write1 <= '1';

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i:
					  waddress <= data_out;
					  data_in <= RR;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);
					  write1 <= '1';

				 END IF;
				state := exec2;
			END IF;
			
--========================================================================
-- MOV
--========================================================================         
			IF (IR(7 DOWNTO 4) = MOV) THEN

				 IF (IR(3 DOWNTO 0) = "0011") THEN  -- A i: Move o valor imediato para RA
					  RA <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i: Move o valor imediato para RB
					  RB <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i: Move o valor imediato para RR
					  RR <= data_out;
					  PC <= STD_LOGIC_VECTOR(unsigned(PC) + 1);

				 END IF;

				 state := fetch;
			END IF;
			
-- XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX
			
		
	


	
--************************************************************************
-- EXECUTE2 STATE
--************************************************************************								
					
			when exec2 =>
	
			LED1	<= '0';
			LED2	<= '0';
			LED3	<= '0';
			LED4	<= '0';
			LED5	<= '1';
			
--========================================================================
-- LOAD
--========================================================================            
			IF (IR(7 DOWNTO 4) = LOAD) THEN
				  
				 IF (IR(3 DOWNTO 0) = "0011") THEN  -- A i: Carrega para o registrador RA o valor do endereço imediato
					  RA <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "0111") THEN  -- B i: Carrega para o registrador RB o valor do endereço imediato
					  RB <= data_out;

				 ELSIF (IR(3 DOWNTO 0) = "1011") THEN  -- R i: Carrega para o registrador RR o valor do endereço imediato
					  RR <= data_out;

				 END IF;
				state := fetch;
			END IF;

--========================================================================
-- STORE
--========================================================================            
			IF (IR(7 DOWNTO 4) = STORE) THEN
				write1 <= '0';
				state := fetch;
			END IF;
			
-- XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX

END CASE;

END IF;

END PROCESS;
	
--************************************************************************
-- ULA 
--************************************************************************
		PROCESS (X, Y, reset)
			
			VARIABLE AUX : STD_LOGIC_VECTOR(7 downto 0);
			VARIABLE RESULT15 : STD_LOGIC_VECTOR(15 downto 0) := (others => '0');
			VARIABLE SUPERIOR : STD_LOGIC_VECTOR(15 downto 0) := "0000000001111111";
			VARIABLE INFERIOR : STD_LOGIC_VECTOR(15 downto 0) := "1111111100000001";
			VARIABLE X_SOMA : STD_LOGIC_VECTOR(15 downto 0) := "00000000" & X;
			VARIABLE Y_SOMA : STD_LOGIC_VECTOR(15 downto 0) := "00000000" & Y;
			
		BEGIN
		
		IF(reset = '1') THEN

			FRover  <= '0';
			FRzero  <= '0';
			FRmaior <= '0';
			FRmenor <= '0';

		END IF;
--========================================================================
-- ARITH 
--========================================================================
			IF(INIT_ULA = '1') THEN
				IF(IR(7 DOWNTO 4) = ADD) THEN
					RESULT15 := STD_LOGIC_VECTOR(signed(X_SOMA) + signed(Y_SOMA));

					-- Trunca RESULT15 para 8 bits e atribui a AUX
					AUX := RESULT15(7 downto 0);

					-- Verificação de overflow usando comparação
					if (signed(RESULT15) > signed(SUPERIOR)) THEN  -- Limite máximo
						FRover <= '1';  -- Overflow: resultado maior que o maior valor positivo
					elsif (signed(RESULT15) < signed(INFERIOR)) THEN  -- Limite mínimo
						FRover <= '1';  -- Overflow: resultado menor que o maior valor negativo
					else
						FRover <= '0';  -- Sem overflow
					end if;
					
					RESULT <= AUX;
					
				ELSIF(IR(7 DOWNTO 4) = SUB or IR(7 DOWNTO 4) = CMP) THEN
					RESULT15 := STD_LOGIC_VECTOR(signed(X_SOMA) - signed(Y_SOMA));
					
					if (signed(RESULT15) > signed(SUPERIOR)) THEN  -- Limite máximo
						FRover <= '1';  -- Overflow: resultado maior que o maior valor positivo
					elsif (signed(RESULT15) < signed(INFERIOR)) THEN  -- Limite mínimo
						FRover <= '1';  -- Overflow: resultado menor que o maior valor negativo
					else
						FRover <= '0';  -- Sem overflow
					end if;
					
					--saidaRR <= RESULT15(7 downto 0);
					--saidaA <= RESULT15(15 downto 8);
					
					if (RESULT15(15) = '1') then
						FRzero <= '0';
						FRmaior <= '0';
						FRmenor <= '1';
						AUX := STD_LOGIC_VECTOR(unsigned(NOT RESULT15(7 downto 0))+1);
					elsif (RESULT15(15 DOWNTO 0) = "0000000000000000") then
						FRzero <= '1';
						FRmaior <= '0';
						FRmenor <= '0';
						AUX := STD_LOGIC_VECTOR(RESULT15(7 downto 0));
					else
						FRzero <= '0';
						FRmaior <= '1';
						FRmenor <= '0';
						AUX := STD_LOGIC_VECTOR(RESULT15(7 downto 0));
					end if;
					
					RESULT <= AUX;
					
				ELSIF(IR(7 DOWNTO 4) = AND1) THEN
				
					RESULT <= X AND Y;
					
				ELSIF(IR(7 DOWNTO 4) = OR1) THEN
				
					RESULT <= X OR Y;
				
				ELSIF(IR(7 DOWNTO 4) = NOT1) THEN
				
					RESULT <= NOT X;

				END IF;
					--saidaRR <= RESULT;
			ELSE
					--saidaRR <= RR;
			END IF;
END PROCESS;
	saidaRR <= RR;
	saidaA <= RA;
	zero <= FRzero;
	maior <= FRmaior;
	menor <= FRmenor;
	over <= FRover;

end main;